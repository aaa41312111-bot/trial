package my_pkg;
    `include "reg_item.v"
    `include "monitor.v"
    `include "driver.v"
    `include "generator.v"
    `include "scoreboard.v"
    `include "env.v"
    `include "something.sv"
endpackage
